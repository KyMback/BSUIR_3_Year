-- megafunction wizard: %ALTECC%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altecc_encoder 

-- ============================================================
-- File Name: altecc_encoder0.vhd
-- Megafunction Name(s):
-- 			altecc_encoder
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 222 10/21/2009 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altecc_encoder CBX_AUTO_BLACKBOX="ALL" device_family="Stratix" lpm_pipeline=0 width_codeword=6 width_dataword=2 data q
--VERSION_BEGIN 9.1 cbx_altecc_encoder 2009:10:21:21:22:16:SJ cbx_mgl 2009:10:21:21:37:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altecc_encoder0_altecc_encoder_31b IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END altecc_encoder0_altecc_encoder_31b;

 ARCHITECTURE RTL OF altecc_encoder0_altecc_encoder_31b IS

	 SIGNAL  wire_w_lg_w_data_wire_range6w8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_q_wire_range19w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_q_wire_range9w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_q_wire_range12w25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_q_wire_range15w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  parity_01_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  parity_02_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  parity_03_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  parity_final_wire :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  q_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_data_wire_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_parity_01_wire_range4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_parity_final_wire_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_parity_final_wire_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_parity_final_wire_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_parity_final_wire_range24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_q_wire_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_q_wire_range9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_q_wire_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_q_wire_range15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_w_lg_w_data_wire_range6w8w(0) <= wire_w_data_wire_range6w(0) XOR wire_w_parity_01_wire_range4w(0);
	wire_w_lg_w_q_wire_range19w21w(0) <= wire_w_q_wire_range19w(0) XOR wire_w_parity_final_wire_range17w(0);
	wire_w_lg_w_q_wire_range9w23w(0) <= wire_w_q_wire_range9w(0) XOR wire_w_parity_final_wire_range20w(0);
	wire_w_lg_w_q_wire_range12w25w(0) <= wire_w_q_wire_range12w(0) XOR wire_w_parity_final_wire_range22w(0);
	wire_w_lg_w_q_wire_range15w27w(0) <= wire_w_q_wire_range15w(0) XOR wire_w_parity_final_wire_range24w(0);
	data_wire <= data;
	parity_01_wire <= ( wire_w_lg_w_data_wire_range6w8w & data_wire(0));
	parity_02_wire(0) <= ( data_wire(0));
	parity_03_wire(0) <= ( data_wire(1));
	parity_final_wire <= ( wire_w_lg_w_q_wire_range15w27w & wire_w_lg_w_q_wire_range12w25w & wire_w_lg_w_q_wire_range9w23w & wire_w_lg_w_q_wire_range19w21w & q_wire(0));
	q <= q_wire;
	q_wire <= ( parity_final_wire(4) & parity_03_wire(0) & parity_02_wire(0) & parity_01_wire(1) & data_wire);
	wire_w_data_wire_range6w(0) <= data_wire(1);
	wire_w_parity_01_wire_range4w(0) <= parity_01_wire(0);
	wire_w_parity_final_wire_range17w(0) <= parity_final_wire(0);
	wire_w_parity_final_wire_range20w(0) <= parity_final_wire(1);
	wire_w_parity_final_wire_range22w(0) <= parity_final_wire(2);
	wire_w_parity_final_wire_range24w(0) <= parity_final_wire(3);
	wire_w_q_wire_range19w(0) <= q_wire(1);
	wire_w_q_wire_range9w(0) <= q_wire(2);
	wire_w_q_wire_range12w(0) <= q_wire(3);
	wire_w_q_wire_range15w(0) <= q_wire(4);

 END RTL; --altecc_encoder0_altecc_encoder_31b
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altecc_encoder0 IS
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		q		: OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
	);
END altecc_encoder0;


ARCHITECTURE RTL OF altecc_encoder0 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (5 DOWNTO 0);



	COMPONENT altecc_encoder0_altecc_encoder_31b
	PORT (
			q	: OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
			data	: IN STD_LOGIC_VECTOR (1 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	q    <= sub_wire0(5 DOWNTO 0);

	altecc_encoder0_altecc_encoder_31b_component : altecc_encoder0_altecc_encoder_31b
	PORT MAP (
		data => data,
		q => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: CONSTANT: lpm_pipeline NUMERIC "0"
-- Retrieval info: CONSTANT: width_codeword NUMERIC "6"
-- Retrieval info: CONSTANT: width_dataword NUMERIC "2"
-- Retrieval info: USED_PORT: data 0 0 2 0 INPUT NODEFVAL "data[1..0]"
-- Retrieval info: USED_PORT: q 0 0 6 0 OUTPUT NODEFVAL "q[5..0]"
-- Retrieval info: CONNECT: @data 0 0 2 0 data 0 0 2 0
-- Retrieval info: CONNECT: q 0 0 6 0 @q 0 0 6 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altecc_encoder0.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altecc_encoder0.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altecc_encoder0.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altecc_encoder0.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altecc_encoder0_inst.vhd FALSE
